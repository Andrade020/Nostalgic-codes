library verilog;
use verilog.vl_types.all;
entity Proc_Simples_vlg_vec_tst is
end Proc_Simples_vlg_vec_tst;
